.title KiCad schematic
M1 /X /A /VDD /VDD PMOS l=1u w=6u
M2 /X /A /VSS /VSS NMOS l=1u w=2u
.end
