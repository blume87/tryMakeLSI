*

.subckt Inv
+       A ; input
+       VDD ; input
+       VSS ; input
+       X ; output


M1 X A VDD VDD PMOS_OR1 l=1u w=6u
M2 X A VSS VSS NMOS_OR1 l=1u w=2u

.ends
